// MKRVIDOR4000_graphics_lite_sys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module MKRVIDOR4000_graphics_lite_sys (
		input  wire        arb_fb_clk,        //     arb_fb.clk
		input  wire        arb_fb_rdy,        //           .rdy
		output wire [30:0] arb_fb_data,       //           .data
		output wire        arb_fb_dv,         //           .dv
		output wire        arb_fb_start,      //           .start
		input  wire        arb_mipi_clk,      //   arb_mipi.clk
		input  wire [14:0] arb_mipi_data,     //           .data
		input  wire        arb_mipi_dv,       //           .dv
		input  wire        arb_mipi_start,    //           .start
		input  wire        clk_clk,           //        clk.clk
		input  wire        clk_0_clk,         //      clk_0.clk
		input  wire        csi_i2c_scl_i,     //    csi_i2c.scl_i
		output wire        csi_i2c_scl_o,     //           .scl_o
		output wire        csi_i2c_scl_en,    //           .scl_en
		input  wire        csi_i2c_sda_i,     //           .sda_i
		output wire        csi_i2c_sda_o,     //           .sda_o
		output wire        csi_i2c_sda_en,    //           .sda_en
		input  wire [10:0] encoder_encoder_a, //    encoder.encoder_a
		input  wire [10:0] encoder_encoder_b, //           .encoder_b
		input  wire        fb_st_start,       //      fb_st.start
		input  wire [30:0] fb_st_data,        //           .data
		input  wire        fb_st_dv,          //           .dv
		output wire        fb_st_ready,       //           .ready
		output wire [7:0]  fb_vport_blu,      //   fb_vport.blu
		output wire        fb_vport_de,       //           .de
		output wire [7:0]  fb_vport_grn,      //           .grn
		output wire        fb_vport_hs,       //           .hs
		output wire        fb_vport_vs,       //           .vs
		output wire [7:0]  fb_vport_red,      //           .red
		output wire        flash_spi_MOSI,    //  flash_spi.MOSI
		output wire        flash_spi_SCLK,    //           .SCLK
		input  wire        flash_spi_MISO,    //           .MISO
		output wire        flash_spi_CS,      //           .CS
		input  wire        hdmi_i2c_scl_i,    //   hdmi_i2c.scl_i
		output wire        hdmi_i2c_scl_o,    //           .scl_o
		output wire        hdmi_i2c_scl_en,   //           .scl_en
		input  wire        hdmi_i2c_sda_i,    //           .sda_i
		output wire        hdmi_i2c_sda_o,    //           .sda_o
		output wire        hdmi_i2c_sda_en,   //           .sda_en
		input  wire [1:0]  irq_in_port,       //        irq.in_port
		output wire [1:0]  irq_out_port,      //           .out_port
		output wire        mb_ak,             //         mb.ak
		input  wire        mb_rq,             //           .rq
		input  wire        mipi_rx_clk,       //    mipi_rx.clk
		input  wire [1:0]  mipi_rx_data,      //           .data
		output wire [23:0] mipi_st_data,      //    mipi_st.data
		output wire        mipi_st_start,     //           .start
		output wire        mipi_st_dv,        //           .dv
		output wire [11:0] neopixel_data,     //   neopixel.data
		output wire        neopixel_clock,    //           .clock
		output wire        nina_spi_MOSI,     //   nina_spi.MOSI
		output wire        nina_spi_SCLK,     //           .SCLK
		input  wire        nina_spi_MISO,     //           .MISO
		output wire        nina_spi_CS,       //           .CS
		input  wire [31:0] pex_pio_in,        //    pex_pio.in
		output wire [31:0] pex_pio_dir,       //           .dir
		output wire [31:0] pex_pio_out,       //           .out
		output wire [63:0] pex_pio_msel,      //           .msel
		input  wire [23:0] qr_vid_in_data,    //  qr_vid_in.data
		input  wire        qr_vid_in_dv,      //           .dv
		input  wire        qr_vid_in_start,   //           .start
		input  wire        qr_vid_in_reset,   //           .reset
		input  wire        qr_vid_in_clk,     //           .clk
		output wire [23:0] qr_vid_out_data,   // qr_vid_out.data
		output wire        qr_vid_out_dv,     //           .dv
		output wire        qr_vid_out_start,  //           .start
		output wire        qspi_dclk,         //       qspi.dclk
		output wire        qspi_ncs,          //           .ncs
		output wire        qspi_oe,           //           .oe
		output wire [3:0]  qspi_dataout,      //           .dataout
		output wire [3:0]  qspi_dataoe,       //           .dataoe
		input  wire [3:0]  qspi_datain,       //           .datain
		input  wire        reset_reset_n,     //      reset.reset_n
		input  wire        reset_0_reset_n,   //    reset_0.reset_n
		input  wire [31:0] sam_pio_in,        //    sam_pio.in
		output wire [31:0] sam_pio_dir,       //           .dir
		output wire [31:0] sam_pio_out,       //           .out
		output wire [63:0] sam_pio_msel,      //           .msel
		output wire [23:0] sam_pwm_pwm,       //    sam_pwm.pwm
		output wire [11:0] sdram_addr,        //      sdram.addr
		output wire [1:0]  sdram_ba,          //           .ba
		output wire        sdram_cas_n,       //           .cas_n
		output wire        sdram_cke,         //           .cke
		output wire        sdram_cs_n,        //           .cs_n
		inout  wire [15:0] sdram_dq,          //           .dq
		output wire [1:0]  sdram_dqm,         //           .dqm
		output wire        sdram_ras_n,       //           .ras_n
		output wire        sdram_we_n,        //           .we_n
		input  wire        vid_clk,           //        vid.clk
		input  wire [31:0] wm_pio_in,         //     wm_pio.in
		output wire [31:0] wm_pio_dir,        //           .dir
		output wire [31:0] wm_pio_out,        //           .out
		output wire [63:0] wm_pio_msel        //           .msel
	);

	wire  [31:0] jtag_bridge_avalon_master_readdata;                         // mm_interconnect_0:JTAG_BRIDGE_avalon_master_readdata -> JTAG_BRIDGE:iREAD_DATA
	wire         jtag_bridge_avalon_master_waitrequest;                      // mm_interconnect_0:JTAG_BRIDGE_avalon_master_waitrequest -> JTAG_BRIDGE:iWAIT_REQUEST
	wire  [31:0] jtag_bridge_avalon_master_address;                          // JTAG_BRIDGE:oADDRESS -> mm_interconnect_0:JTAG_BRIDGE_avalon_master_address
	wire         jtag_bridge_avalon_master_read;                             // JTAG_BRIDGE:oREAD -> mm_interconnect_0:JTAG_BRIDGE_avalon_master_read
	wire         jtag_bridge_avalon_master_readdatavalid;                    // mm_interconnect_0:JTAG_BRIDGE_avalon_master_readdatavalid -> JTAG_BRIDGE:iREAD_DATA_VALID
	wire         jtag_bridge_avalon_master_write;                            // JTAG_BRIDGE:oWRITE -> mm_interconnect_0:JTAG_BRIDGE_avalon_master_write
	wire  [31:0] jtag_bridge_avalon_master_writedata;                        // JTAG_BRIDGE:oWRITE_DATA -> mm_interconnect_0:JTAG_BRIDGE_avalon_master_writedata
	wire  [31:0] mm_interconnect_0_mb_mst_readdata;                          // mb:oMST_READ_DATA -> mm_interconnect_0:mb_mst_readdata
	wire   [8:0] mm_interconnect_0_mb_mst_address;                           // mm_interconnect_0:mb_mst_address -> mb:iMST_ADDRESS
	wire         mm_interconnect_0_mb_mst_read;                              // mm_interconnect_0:mb_mst_read -> mb:iMST_READ
	wire         mm_interconnect_0_mb_mst_write;                             // mm_interconnect_0:mb_mst_write -> mb:iMST_WRITE
	wire  [31:0] mm_interconnect_0_mb_mst_writedata;                         // mm_interconnect_0:mb_mst_writedata -> mb:iMST_WRITE_DATA
	wire         neopixel_0_data_waitrequest;                                // mm_interconnect_1:NEOPIXEL_0_data_waitrequest -> NEOPIXEL_0:iDATA_WAIT_REQUEST
	wire  [31:0] neopixel_0_data_readdata;                                   // mm_interconnect_1:NEOPIXEL_0_data_readdata -> NEOPIXEL_0:iDATA_READ_DATA
	wire  [31:0] neopixel_0_data_address;                                    // NEOPIXEL_0:oDATA_ADDRESS -> mm_interconnect_1:NEOPIXEL_0_data_address
	wire         neopixel_0_data_read;                                       // NEOPIXEL_0:oDATA_READ -> mm_interconnect_1:NEOPIXEL_0_data_read
	wire         neopixel_0_data_readdatavalid;                              // mm_interconnect_1:NEOPIXEL_0_data_readdatavalid -> NEOPIXEL_0:iDATA_READ_DATA_VALID
	wire   [4:0] neopixel_0_data_burstcount;                                 // NEOPIXEL_0:oDATA_BURST_COUNT -> mm_interconnect_1:NEOPIXEL_0_data_burstcount
	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_1:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_1:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_0_data_master_debugaccess
	wire  [23:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_1:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_1:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_1:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_1:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_1:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_1:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_1:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [23:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_1:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_1:nios2_gen2_0_instruction_master_read
	wire  [15:0] mm_interconnect_1_sdram_arbiter_avl_readdata;               // SDRAM_ARBITER:oAVL_READ_DATA -> mm_interconnect_1:SDRAM_ARBITER_avl_readdata
	wire         mm_interconnect_1_sdram_arbiter_avl_waitrequest;            // SDRAM_ARBITER:oAVL_WAIT_REQUEST -> mm_interconnect_1:SDRAM_ARBITER_avl_waitrequest
	wire  [21:0] mm_interconnect_1_sdram_arbiter_avl_address;                // mm_interconnect_1:SDRAM_ARBITER_avl_address -> SDRAM_ARBITER:iAVL_ADDRESS
	wire         mm_interconnect_1_sdram_arbiter_avl_read;                   // mm_interconnect_1:SDRAM_ARBITER_avl_read -> SDRAM_ARBITER:iAVL_READ
	wire   [1:0] mm_interconnect_1_sdram_arbiter_avl_byteenable;             // mm_interconnect_1:SDRAM_ARBITER_avl_byteenable -> SDRAM_ARBITER:iAVL_BYTE_ENABLE
	wire         mm_interconnect_1_sdram_arbiter_avl_readdatavalid;          // SDRAM_ARBITER:oAVL_READ_DATA_VALID -> mm_interconnect_1:SDRAM_ARBITER_avl_readdatavalid
	wire         mm_interconnect_1_sdram_arbiter_avl_write;                  // mm_interconnect_1:SDRAM_ARBITER_avl_write -> SDRAM_ARBITER:iAVL_WRITE
	wire  [15:0] mm_interconnect_1_sdram_arbiter_avl_writedata;              // mm_interconnect_1:SDRAM_ARBITER_avl_writedata -> SDRAM_ARBITER:iAVL_WRITE_DATA
	wire   [5:0] mm_interconnect_1_sdram_arbiter_avl_burstcount;             // mm_interconnect_1:SDRAM_ARBITER_avl_burstcount -> SDRAM_ARBITER:iAVL_BURST_COUNT
	wire         mm_interconnect_1_csi_i2c_avalon_slave_0_chipselect;        // mm_interconnect_1:csi_i2c_avalon_slave_0_chipselect -> csi_i2c:wb_stb_i
	wire  [31:0] mm_interconnect_1_csi_i2c_avalon_slave_0_readdata;          // csi_i2c:wb_dat_o -> mm_interconnect_1:csi_i2c_avalon_slave_0_readdata
	wire         mm_interconnect_1_csi_i2c_avalon_slave_0_waitrequest;       // csi_i2c:wb_ack_o -> mm_interconnect_1:csi_i2c_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_1_csi_i2c_avalon_slave_0_address;           // mm_interconnect_1:csi_i2c_avalon_slave_0_address -> csi_i2c:wb_adr_i
	wire         mm_interconnect_1_csi_i2c_avalon_slave_0_write;             // mm_interconnect_1:csi_i2c_avalon_slave_0_write -> csi_i2c:wb_we_i
	wire  [31:0] mm_interconnect_1_csi_i2c_avalon_slave_0_writedata;         // mm_interconnect_1:csi_i2c_avalon_slave_0_writedata -> csi_i2c:wb_dat_i
	wire   [4:0] mm_interconnect_1_sam_pwm_avalon_slave_0_address;           // mm_interconnect_1:sam_pwm_avalon_slave_0_address -> sam_pwm:iADDRESS
	wire         mm_interconnect_1_sam_pwm_avalon_slave_0_write;             // mm_interconnect_1:sam_pwm_avalon_slave_0_write -> sam_pwm:iWRITE
	wire  [31:0] mm_interconnect_1_sam_pwm_avalon_slave_0_writedata;         // mm_interconnect_1:sam_pwm_avalon_slave_0_writedata -> sam_pwm:iWRITE_DATA
	wire         mm_interconnect_1_hdmi_i2c_avalon_slave_0_chipselect;       // mm_interconnect_1:hdmi_i2c_avalon_slave_0_chipselect -> hdmi_i2c:wb_stb_i
	wire  [31:0] mm_interconnect_1_hdmi_i2c_avalon_slave_0_readdata;         // hdmi_i2c:wb_dat_o -> mm_interconnect_1:hdmi_i2c_avalon_slave_0_readdata
	wire         mm_interconnect_1_hdmi_i2c_avalon_slave_0_waitrequest;      // hdmi_i2c:wb_ack_o -> mm_interconnect_1:hdmi_i2c_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_1_hdmi_i2c_avalon_slave_0_address;          // mm_interconnect_1:hdmi_i2c_avalon_slave_0_address -> hdmi_i2c:wb_adr_i
	wire         mm_interconnect_1_hdmi_i2c_avalon_slave_0_write;            // mm_interconnect_1:hdmi_i2c_avalon_slave_0_write -> hdmi_i2c:wb_we_i
	wire  [31:0] mm_interconnect_1_hdmi_i2c_avalon_slave_0_writedata;        // mm_interconnect_1:hdmi_i2c_avalon_slave_0_writedata -> hdmi_i2c:wb_dat_i
	wire  [31:0] mm_interconnect_1_quad_encoder_0_avalon_slave_0_readdata;   // QUAD_ENCODER_0:oAVL_READ_DATA -> mm_interconnect_1:QUAD_ENCODER_0_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_1_quad_encoder_0_avalon_slave_0_address;    // mm_interconnect_1:QUAD_ENCODER_0_avalon_slave_0_address -> QUAD_ENCODER_0:iAVL_ADDRESS
	wire         mm_interconnect_1_quad_encoder_0_avalon_slave_0_read;       // mm_interconnect_1:QUAD_ENCODER_0_avalon_slave_0_read -> QUAD_ENCODER_0:iAVL_READ
	wire  [31:0] mm_interconnect_1_qspi_avl_csr_readdata;                    // qspi:avl_csr_rddata -> mm_interconnect_1:qspi_avl_csr_readdata
	wire         mm_interconnect_1_qspi_avl_csr_waitrequest;                 // qspi:avl_csr_waitrequest -> mm_interconnect_1:qspi_avl_csr_waitrequest
	wire   [3:0] mm_interconnect_1_qspi_avl_csr_address;                     // mm_interconnect_1:qspi_avl_csr_address -> qspi:avl_csr_addr
	wire         mm_interconnect_1_qspi_avl_csr_read;                        // mm_interconnect_1:qspi_avl_csr_read -> qspi:avl_csr_read
	wire         mm_interconnect_1_qspi_avl_csr_readdatavalid;               // qspi:avl_csr_rddata_valid -> mm_interconnect_1:qspi_avl_csr_readdatavalid
	wire         mm_interconnect_1_qspi_avl_csr_write;                       // mm_interconnect_1:qspi_avl_csr_write -> qspi:avl_csr_write
	wire  [31:0] mm_interconnect_1_qspi_avl_csr_writedata;                   // mm_interconnect_1:qspi_avl_csr_writedata -> qspi:avl_csr_wrdata
	wire  [31:0] mm_interconnect_1_qspi_avl_mem_readdata;                    // qspi:avl_mem_rddata -> mm_interconnect_1:qspi_avl_mem_readdata
	wire         mm_interconnect_1_qspi_avl_mem_waitrequest;                 // qspi:avl_mem_waitrequest -> mm_interconnect_1:qspi_avl_mem_waitrequest
	wire  [18:0] mm_interconnect_1_qspi_avl_mem_address;                     // mm_interconnect_1:qspi_avl_mem_address -> qspi:avl_mem_addr
	wire         mm_interconnect_1_qspi_avl_mem_read;                        // mm_interconnect_1:qspi_avl_mem_read -> qspi:avl_mem_read
	wire   [3:0] mm_interconnect_1_qspi_avl_mem_byteenable;                  // mm_interconnect_1:qspi_avl_mem_byteenable -> qspi:avl_mem_byteenable
	wire         mm_interconnect_1_qspi_avl_mem_readdatavalid;               // qspi:avl_mem_rddata_valid -> mm_interconnect_1:qspi_avl_mem_readdatavalid
	wire         mm_interconnect_1_qspi_avl_mem_write;                       // mm_interconnect_1:qspi_avl_mem_write -> qspi:avl_mem_write
	wire  [31:0] mm_interconnect_1_qspi_avl_mem_writedata;                   // mm_interconnect_1:qspi_avl_mem_writedata -> qspi:avl_mem_wrdata
	wire   [6:0] mm_interconnect_1_qspi_avl_mem_burstcount;                  // mm_interconnect_1:qspi_avl_mem_burstcount -> qspi:avl_mem_burstcount
	wire  [31:0] mm_interconnect_1_sysid_qsys_0_control_slave_readdata;      // sysid_qsys_0:readdata -> mm_interconnect_1:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_qsys_0_control_slave_address;       // mm_interconnect_1:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_1_neopixel_0_csr_readdata;                  // NEOPIXEL_0:oCSR_READ_DATA -> mm_interconnect_1:NEOPIXEL_0_csr_readdata
	wire   [3:0] mm_interconnect_1_neopixel_0_csr_address;                   // mm_interconnect_1:NEOPIXEL_0_csr_address -> NEOPIXEL_0:iCSR_ADDRESS
	wire         mm_interconnect_1_neopixel_0_csr_read;                      // mm_interconnect_1:NEOPIXEL_0_csr_read -> NEOPIXEL_0:iCSR_READ
	wire         mm_interconnect_1_neopixel_0_csr_write;                     // mm_interconnect_1:NEOPIXEL_0_csr_write -> NEOPIXEL_0:iCSR_WRITE
	wire  [31:0] mm_interconnect_1_neopixel_0_csr_writedata;                 // mm_interconnect_1:NEOPIXEL_0_csr_writedata -> NEOPIXEL_0:iCSR_WRITE_DATA
	wire  [31:0] mm_interconnect_1_qrcode_finder_0_ctrl_readdata;            // QRCODE_FINDER_0:oREAD_DATA -> mm_interconnect_1:QRCODE_FINDER_0_ctrl_readdata
	wire  [10:0] mm_interconnect_1_qrcode_finder_0_ctrl_address;             // mm_interconnect_1:QRCODE_FINDER_0_ctrl_address -> QRCODE_FINDER_0:iADDRESS
	wire         mm_interconnect_1_qrcode_finder_0_ctrl_read;                // mm_interconnect_1:QRCODE_FINDER_0_ctrl_read -> QRCODE_FINDER_0:iREAD
	wire         mm_interconnect_1_qrcode_finder_0_ctrl_write;               // mm_interconnect_1:QRCODE_FINDER_0_ctrl_write -> QRCODE_FINDER_0:iWRITE
	wire  [31:0] mm_interconnect_1_qrcode_finder_0_ctrl_writedata;           // mm_interconnect_1:QRCODE_FINDER_0_ctrl_writedata -> QRCODE_FINDER_0:iWRITE_DATA
	wire         mm_interconnect_1_nina_spi_d_chipselect;                    // mm_interconnect_1:nina_spi_d_chipselect -> nina_spi:stb_i
	wire  [31:0] mm_interconnect_1_nina_spi_d_readdata;                      // nina_spi:dat_o -> mm_interconnect_1:nina_spi_d_readdata
	wire   [2:0] mm_interconnect_1_nina_spi_d_address;                       // mm_interconnect_1:nina_spi_d_address -> nina_spi:adr_i
	wire         mm_interconnect_1_nina_spi_d_write;                         // mm_interconnect_1:nina_spi_d_write -> nina_spi:we_i
	wire  [31:0] mm_interconnect_1_nina_spi_d_writedata;                     // mm_interconnect_1:nina_spi_d_writedata -> nina_spi:dat_i
	wire         mm_interconnect_1_flash_spi_d_chipselect;                   // mm_interconnect_1:flash_spi_d_chipselect -> flash_spi:stb_i
	wire  [31:0] mm_interconnect_1_flash_spi_d_readdata;                     // flash_spi:dat_o -> mm_interconnect_1:flash_spi_d_readdata
	wire   [2:0] mm_interconnect_1_flash_spi_d_address;                      // mm_interconnect_1:flash_spi_d_address -> flash_spi:adr_i
	wire         mm_interconnect_1_flash_spi_d_write;                        // mm_interconnect_1:flash_spi_d_write -> flash_spi:we_i
	wire  [31:0] mm_interconnect_1_flash_spi_d_writedata;                    // mm_interconnect_1:flash_spi_d_writedata -> flash_spi:dat_i
	wire  [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_1_sam_pio_s1_readdata;                      // sam_pio:oREAD_DATA -> mm_interconnect_1:sam_pio_s1_readdata
	wire   [2:0] mm_interconnect_1_sam_pio_s1_address;                       // mm_interconnect_1:sam_pio_s1_address -> sam_pio:iADDRESS
	wire         mm_interconnect_1_sam_pio_s1_read;                          // mm_interconnect_1:sam_pio_s1_read -> sam_pio:iREAD
	wire         mm_interconnect_1_sam_pio_s1_write;                         // mm_interconnect_1:sam_pio_s1_write -> sam_pio:iWRITE
	wire  [31:0] mm_interconnect_1_sam_pio_s1_writedata;                     // mm_interconnect_1:sam_pio_s1_writedata -> sam_pio:iWRITE_DATA
	wire  [31:0] mm_interconnect_1_pex_pio_s1_readdata;                      // pex_pio:oREAD_DATA -> mm_interconnect_1:pex_pio_s1_readdata
	wire   [2:0] mm_interconnect_1_pex_pio_s1_address;                       // mm_interconnect_1:pex_pio_s1_address -> pex_pio:iADDRESS
	wire         mm_interconnect_1_pex_pio_s1_read;                          // mm_interconnect_1:pex_pio_s1_read -> pex_pio:iREAD
	wire         mm_interconnect_1_pex_pio_s1_write;                         // mm_interconnect_1:pex_pio_s1_write -> pex_pio:iWRITE
	wire  [31:0] mm_interconnect_1_pex_pio_s1_writedata;                     // mm_interconnect_1:pex_pio_s1_writedata -> pex_pio:iWRITE_DATA
	wire  [31:0] mm_interconnect_1_wm_pio_s1_readdata;                       // wm_pio:oREAD_DATA -> mm_interconnect_1:wm_pio_s1_readdata
	wire   [2:0] mm_interconnect_1_wm_pio_s1_address;                        // mm_interconnect_1:wm_pio_s1_address -> wm_pio:iADDRESS
	wire         mm_interconnect_1_wm_pio_s1_read;                           // mm_interconnect_1:wm_pio_s1_read -> wm_pio:iREAD
	wire         mm_interconnect_1_wm_pio_s1_write;                          // mm_interconnect_1:wm_pio_s1_write -> wm_pio:iWRITE
	wire  [31:0] mm_interconnect_1_wm_pio_s1_writedata;                      // mm_interconnect_1:wm_pio_s1_writedata -> wm_pio:iWRITE_DATA
	wire         mm_interconnect_1_irq_s1_chipselect;                        // mm_interconnect_1:irq_s1_chipselect -> irq:chipselect
	wire  [31:0] mm_interconnect_1_irq_s1_readdata;                          // irq:readdata -> mm_interconnect_1:irq_s1_readdata
	wire   [1:0] mm_interconnect_1_irq_s1_address;                           // mm_interconnect_1:irq_s1_address -> irq:address
	wire         mm_interconnect_1_irq_s1_write;                             // mm_interconnect_1:irq_s1_write -> irq:write_n
	wire  [31:0] mm_interconnect_1_irq_s1_writedata;                         // mm_interconnect_1:irq_s1_writedata -> irq:writedata
	wire         mm_interconnect_1_onchip_memory2_0_s1_chipselect;           // mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_readdata;             // onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_1_onchip_memory2_0_s1_address;              // mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_1_onchip_memory2_0_s1_byteenable;           // mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_1_onchip_memory2_0_s1_write;                // mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_writedata;            // mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_1_onchip_memory2_0_s1_clken;                // mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_1_timer_0_s1_chipselect;                    // mm_interconnect_1:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_1_timer_0_s1_readdata;                      // timer_0:readdata -> mm_interconnect_1:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_0_s1_address;                       // mm_interconnect_1:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_1_timer_0_s1_write;                         // mm_interconnect_1:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_1_timer_0_s1_writedata;                     // mm_interconnect_1:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] mm_interconnect_1_mb_slv_readdata;                          // mb:oSLV_READ_DATA -> mm_interconnect_1:mb_slv_readdata
	wire   [8:0] mm_interconnect_1_mb_slv_address;                           // mm_interconnect_1:mb_slv_address -> mb:iSLV_ADDRESS
	wire         mm_interconnect_1_mb_slv_read;                              // mm_interconnect_1:mb_slv_read -> mb:iSLV_READ
	wire         mm_interconnect_1_mb_slv_write;                             // mm_interconnect_1:mb_slv_write -> mb:iSLV_WRITE
	wire  [31:0] mm_interconnect_1_mb_slv_writedata;                         // mm_interconnect_1:mb_slv_writedata -> mb:iSLV_WRITE_DATA
	wire         mm_interconnect_1_onchip_memory2_0_s2_chipselect;           // mm_interconnect_1:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s2_readdata;             // onchip_memory2_0:readdata2 -> mm_interconnect_1:onchip_memory2_0_s2_readdata
	wire  [11:0] mm_interconnect_1_onchip_memory2_0_s2_address;              // mm_interconnect_1:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	wire   [3:0] mm_interconnect_1_onchip_memory2_0_s2_byteenable;           // mm_interconnect_1:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	wire         mm_interconnect_1_onchip_memory2_0_s2_write;                // mm_interconnect_1:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s2_writedata;            // mm_interconnect_1:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	wire         mm_interconnect_1_onchip_memory2_0_s2_clken;                // mm_interconnect_1:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	wire  [15:0] sdram_arbiter_sdram_readdata;                               // mm_interconnect_2:SDRAM_ARBITER_sdram_readdata -> SDRAM_ARBITER:iSDRAM_READ_DATA
	wire         sdram_arbiter_sdram_waitrequest;                            // mm_interconnect_2:SDRAM_ARBITER_sdram_waitrequest -> SDRAM_ARBITER:iSDRAM_WAIT_REQUEST
	wire  [21:0] sdram_arbiter_sdram_address;                                // SDRAM_ARBITER:oSDRAM_ADDRESS -> mm_interconnect_2:SDRAM_ARBITER_sdram_address
	wire         sdram_arbiter_sdram_read;                                   // SDRAM_ARBITER:oSDRAM_READ -> mm_interconnect_2:SDRAM_ARBITER_sdram_read
	wire   [1:0] sdram_arbiter_sdram_byteenable;                             // SDRAM_ARBITER:oSDRAM_BYTE_ENABLE -> mm_interconnect_2:SDRAM_ARBITER_sdram_byteenable
	wire         sdram_arbiter_sdram_readdatavalid;                          // mm_interconnect_2:SDRAM_ARBITER_sdram_readdatavalid -> SDRAM_ARBITER:iSDRAM_READ_DATA_VALID
	wire         sdram_arbiter_sdram_write;                                  // SDRAM_ARBITER:oSDRAM_WRITE -> mm_interconnect_2:SDRAM_ARBITER_sdram_write
	wire  [15:0] sdram_arbiter_sdram_writedata;                              // SDRAM_ARBITER:oSDRAM_WRITE_DATA -> mm_interconnect_2:SDRAM_ARBITER_sdram_writedata
	wire         mm_interconnect_2_sdram_s1_chipselect;                      // mm_interconnect_2:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_2_sdram_s1_readdata;                        // sdram:za_data -> mm_interconnect_2:sdram_s1_readdata
	wire         mm_interconnect_2_sdram_s1_waitrequest;                     // sdram:za_waitrequest -> mm_interconnect_2:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_2_sdram_s1_address;                         // mm_interconnect_2:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_2_sdram_s1_read;                            // mm_interconnect_2:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_2_sdram_s1_byteenable;                      // mm_interconnect_2:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_2_sdram_s1_readdatavalid;                   // sdram:za_valid -> mm_interconnect_2:sdram_s1_readdatavalid
	wire         mm_interconnect_2_sdram_s1_write;                           // mm_interconnect_2:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_2_sdram_s1_writedata;                       // mm_interconnect_2:sdram_s1_writedata -> sdram:az_data
	wire         irq_mapper_receiver0_irq;                                   // NEOPIXEL_0:oIRQ -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // irq:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                   // nina_spi:int_o -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                   // timer_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [JTAG_BRIDGE:iRESET, NEOPIXEL_0:iRESET, QRCODE_FINDER_0:iRESET, QUAD_ENCODER_0:iRESET, SDRAM_ARBITER:iRESET, csi_i2c:wb_rst_i, flash_spi:rst_i, hdmi_i2c:wb_rst_i, irq:reset_n, mb:iRESET, mm_interconnect_0:JTAG_BRIDGE_reset_reset_bridge_in_reset_reset, mm_interconnect_1:NEOPIXEL_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:SDRAM_ARBITER_reset_reset_bridge_in_reset_reset, nina_spi:rst_i, onchip_memory2_0:reset, onchip_memory2_0:reset2, pex_pio:iRESET, rst_translator:in_reset, sam_pio:iRESET, sam_pwm:iRESET, sdram:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, wm_pio:iRESET]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_0:reset_req2, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                     // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in1
	wire         rst_controller_002_reset_out_reset;                         // rst_controller_002:reset_out -> [mm_interconnect_1:qspi_reset_reset_bridge_in_reset_reset, qspi:reset_n]

	FBST #(
		.pHRES   (640),
		.pVRES   (480),
		.pHTOTAL (762),
		.pVTOTAL (525),
		.pHSS    (656),
		.pHSE    (752),
		.pVSS    (490),
		.pVSE    (492)
	) fbst_0 (
		.oBLU          (fb_vport_blu), //   vport.blu
		.oDE           (fb_vport_de),  //        .de
		.oGRN          (fb_vport_grn), //        .grn
		.oHS           (fb_vport_hs),  //        .hs
		.oVS           (fb_vport_vs),  //        .vs
		.oRED          (fb_vport_red), //        .red
		.iCLK          (vid_clk),      // vid_clk.clk
		.iFB_START     (fb_st_start),  //  stream.start
		.iFB_DATA      (fb_st_data),   //        .data
		.iFB_DATAVALID (fb_st_dv),     //        .dv
		.oFB_READY     (fb_st_ready)   //        .ready
	);

	JTAG_BRIDGE jtag_bridge (
		.oADDRESS          (jtag_bridge_avalon_master_address),       // avalon_master.address
		.oWRITE            (jtag_bridge_avalon_master_write),         //              .write
		.oREAD             (jtag_bridge_avalon_master_read),          //              .read
		.oWRITE_DATA       (jtag_bridge_avalon_master_writedata),     //              .writedata
		.iREAD_DATA        (jtag_bridge_avalon_master_readdata),      //              .readdata
		.iWAIT_REQUEST     (jtag_bridge_avalon_master_waitrequest),   //              .waitrequest
		.iREAD_DATA_VALID  (jtag_bridge_avalon_master_readdatavalid), //              .readdatavalid
		.iEVENT_WRITE_DATA (),                                        //         event.writedata
		.iEVENT_WRITE      (),                                        //              .write
		.oEVENT_EMPTY      (),                                        //           irq.irq
		.iRESET            (rst_controller_reset_out_reset),          //         reset.reset
		.iCLK              (clk_clk)                                  //         clock.clk
	);

	MIPI_RX mipi_rx_st_0 (
		.iMIPI_CLK        (mipi_rx_clk),   //    mipi.clk
		.iMIPI_D          (mipi_rx_data),  //        .data
		.oMIPI_DATA       (mipi_st_data),  // mipi_st.data
		.oMIPI_START      (mipi_st_start), //        .start
		.oMIPI_DATA_VALID (mipi_st_dv)     //        .dv
	);

	NEOPIXEL #(
		.pCHANNELS      (11),
		.pSTART_ADDRESS (2097152)
	) neopixel_0 (
		.oCSR_READ_DATA        (mm_interconnect_1_neopixel_0_csr_readdata),  //   csr.readdata
		.iCSR_WRITE_DATA       (mm_interconnect_1_neopixel_0_csr_writedata), //      .writedata
		.iCSR_ADDRESS          (mm_interconnect_1_neopixel_0_csr_address),   //      .address
		.iCSR_READ             (mm_interconnect_1_neopixel_0_csr_read),      //      .read
		.iCSR_WRITE            (mm_interconnect_1_neopixel_0_csr_write),     //      .write
		.iCLOCK                (clk_clk),                                    // clock.clk
		.iRESET                (rst_controller_reset_out_reset),             // reset.reset
		.oDATA                 (neopixel_data),                              // pixel.data
		.oCLK                  (neopixel_clock),                             //      .clock
		.oDATA_ADDRESS         (neopixel_0_data_address),                    //  data.address
		.oDATA_READ            (neopixel_0_data_read),                       //      .read
		.iDATA_WAIT_REQUEST    (neopixel_0_data_waitrequest),                //      .waitrequest
		.oDATA_BURST_COUNT     (neopixel_0_data_burstcount),                 //      .burstcount
		.iDATA_READ_DATA       (neopixel_0_data_readdata),                   //      .readdata
		.iDATA_READ_DATA_VALID (neopixel_0_data_readdatavalid),              //      .readdatavalid
		.oIRQ                  (irq_mapper_receiver0_irq)                    //   irq.irq
	);

	QRCODE_FINDER #(
		.pHRES      (640),
		.pVRES      (480),
		.pTHRESHOLD (60)
	) qrcode_finder_0 (
		.iADDRESS        (mm_interconnect_1_qrcode_finder_0_ctrl_address),   //    ctrl.address
		.iWRITE_DATA     (mm_interconnect_1_qrcode_finder_0_ctrl_writedata), //        .writedata
		.iWRITE          (mm_interconnect_1_qrcode_finder_0_ctrl_write),     //        .write
		.iREAD           (mm_interconnect_1_qrcode_finder_0_ctrl_read),      //        .read
		.oREAD_DATA      (mm_interconnect_1_qrcode_finder_0_ctrl_readdata),  //        .readdata
		.iRESET          (rst_controller_reset_out_reset),                   //   reset.reset
		.iCLOCK          (clk_clk),                                          //   clock.clk
		.iVID_DATA       (qr_vid_in_data),                                   //  vid_in.data
		.iVID_DATA_VALID (qr_vid_in_dv),                                     //        .dv
		.iVID_START      (qr_vid_in_start),                                  //        .start
		.iVID_RESET      (qr_vid_in_reset),                                  //        .reset
		.iVID_CLOCK      (qr_vid_in_clk),                                    //        .clk
		.oVID_DATA       (qr_vid_out_data),                                  // vid_out.data
		.oVID_DATA_VALID (qr_vid_out_dv),                                    //        .dv
		.oVID_START      (qr_vid_out_start)                                  //        .start
	);

	QUAD_ENCODER #(
		.pENCODERS          (11),
		.pENCODER_PRECISION (32)
	) quad_encoder_0 (
		.oAVL_READ_DATA (mm_interconnect_1_quad_encoder_0_avalon_slave_0_readdata), // avalon_slave_0.readdata
		.iAVL_READ      (mm_interconnect_1_quad_encoder_0_avalon_slave_0_read),     //               .read
		.iAVL_ADDRESS   (mm_interconnect_1_quad_encoder_0_avalon_slave_0_address),  //               .address
		.iCLOCK         (clk_clk),                                                  //     clock_sink.clk
		.iRESET         (rst_controller_reset_out_reset),                           //     reset_sink.reset
		.iENCODER_A     (encoder_encoder_a),                                        //        encoder.encoder_a
		.iENCODER_B     (encoder_encoder_b)                                         //               .encoder_b
	);

	SDRAM_ARBITER #(
		.pBURST_SIZE   (128),
		.pCAM_OFFSET_A (0),
		.pCAM_OFFSET_B (307200),
		.pFB_OFFSET    (614400),
		.pFB_SIZE      (307200),
		.pADDRESS_BITS (22)
	) sdram_arbiter (
		.oSDRAM_ADDRESS         (sdram_arbiter_sdram_address),                       // sdram.address
		.oSDRAM_WRITE           (sdram_arbiter_sdram_write),                         //      .write
		.oSDRAM_READ            (sdram_arbiter_sdram_read),                          //      .read
		.oSDRAM_WRITE_DATA      (sdram_arbiter_sdram_writedata),                     //      .writedata
		.iSDRAM_READ_DATA       (sdram_arbiter_sdram_readdata),                      //      .readdata
		.iSDRAM_WAIT_REQUEST    (sdram_arbiter_sdram_waitrequest),                   //      .waitrequest
		.iSDRAM_READ_DATA_VALID (sdram_arbiter_sdram_readdatavalid),                 //      .readdatavalid
		.oSDRAM_BYTE_ENABLE     (sdram_arbiter_sdram_byteenable),                    //      .byteenable
		.iMEM_CLK               (clk_clk),                                           // clock.clk
		.iRESET                 (rst_controller_reset_out_reset),                    // reset.reset
		.iFB_CLK                (arb_fb_clk),                                        //    fb.clk
		.iFB_READY              (arb_fb_rdy),                                        //      .rdy
		.oFB_DATA               (arb_fb_data),                                       //      .data
		.oFB_DATA_VALID         (arb_fb_dv),                                         //      .dv
		.oFB_START              (arb_fb_start),                                      //      .start
		.iMIPI_CLK              (arb_mipi_clk),                                      //  mipi.clk
		.iMIPI_DATA             (arb_mipi_data),                                     //      .data
		.iMIPI_DATA_VALID       (arb_mipi_dv),                                       //      .dv
		.iMIPI_START            (arb_mipi_start),                                    //      .start
		.oAVL_READ_DATA         (mm_interconnect_1_sdram_arbiter_avl_readdata),      //   avl.readdata
		.oAVL_READ_DATA_VALID   (mm_interconnect_1_sdram_arbiter_avl_readdatavalid), //      .readdatavalid
		.iAVL_WRITE_DATA        (mm_interconnect_1_sdram_arbiter_avl_writedata),     //      .writedata
		.oAVL_WAIT_REQUEST      (mm_interconnect_1_sdram_arbiter_avl_waitrequest),   //      .waitrequest
		.iAVL_ADDRESS           (mm_interconnect_1_sdram_arbiter_avl_address),       //      .address
		.iAVL_BURST_COUNT       (mm_interconnect_1_sdram_arbiter_avl_burstcount),    //      .burstcount
		.iAVL_READ              (mm_interconnect_1_sdram_arbiter_avl_read),          //      .read
		.iAVL_WRITE             (mm_interconnect_1_sdram_arbiter_avl_write),         //      .write
		.iAVL_BYTE_ENABLE       (mm_interconnect_1_sdram_arbiter_avl_byteenable)     //      .byteenable
	);

	o_i2c_master csi_i2c (
		.wb_clk_i     (clk_clk),                                              //       clock_sink.clk
		.wb_rst_i     (rst_controller_reset_out_reset),                       // clock_sink_reset.reset
		.wb_ack_o     (mm_interconnect_1_csi_i2c_avalon_slave_0_waitrequest), //   avalon_slave_0.waitrequest_n
		.wb_adr_i     (mm_interconnect_1_csi_i2c_avalon_slave_0_address),     //                 .address
		.wb_dat_i     (mm_interconnect_1_csi_i2c_avalon_slave_0_writedata),   //                 .writedata
		.wb_stb_i     (mm_interconnect_1_csi_i2c_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_we_i      (mm_interconnect_1_csi_i2c_avalon_slave_0_write),       //                 .write
		.wb_dat_o     (mm_interconnect_1_csi_i2c_avalon_slave_0_readdata),    //                 .readdata
		.scl_pad_i    (csi_i2c_scl_i),                                        //    conduit_start.scl_i
		.scl_pad_o    (csi_i2c_scl_o),                                        //                 .scl_o
		.scl_padoen_o (csi_i2c_scl_en),                                       //                 .scl_en
		.sda_pad_i    (csi_i2c_sda_i),                                        //                 .sda_i
		.sda_pad_o    (csi_i2c_sda_o),                                        //                 .sda_o
		.sda_padoen_o (csi_i2c_sda_en),                                       //                 .sda_en
		.wb_inta_o    ()                                                      // interrupt_sender.irq
	);

	tiny_spi #(
		.BAUD_WIDTH (8),
		.BAUD_DIV   (0),
		.SPI_MODE   (0)
	) flash_spi (
		.stb_i (mm_interconnect_1_flash_spi_d_chipselect), //     d.chipselect
		.we_i  (mm_interconnect_1_flash_spi_d_write),      //      .write
		.dat_i (mm_interconnect_1_flash_spi_d_writedata),  //      .writedata
		.adr_i (mm_interconnect_1_flash_spi_d_address),    //      .address
		.dat_o (mm_interconnect_1_flash_spi_d_readdata),   //      .readdata
		.clk_i (clk_clk),                                  //   clk.clk
		.rst_i (rst_controller_reset_out_reset),           // reset.reset
		.int_o (),                                         //   irq.irq
		.MOSI  (flash_spi_MOSI),                           //   spi.MOSI
		.SCLK  (flash_spi_SCLK),                           //      .SCLK
		.MISO  (flash_spi_MISO),                           //      .MISO
		.CS    (flash_spi_CS)                              //      .CS
	);

	o_i2c_master hdmi_i2c (
		.wb_clk_i     (clk_clk),                                               //       clock_sink.clk
		.wb_rst_i     (rst_controller_reset_out_reset),                        // clock_sink_reset.reset
		.wb_ack_o     (mm_interconnect_1_hdmi_i2c_avalon_slave_0_waitrequest), //   avalon_slave_0.waitrequest_n
		.wb_adr_i     (mm_interconnect_1_hdmi_i2c_avalon_slave_0_address),     //                 .address
		.wb_dat_i     (mm_interconnect_1_hdmi_i2c_avalon_slave_0_writedata),   //                 .writedata
		.wb_stb_i     (mm_interconnect_1_hdmi_i2c_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_we_i      (mm_interconnect_1_hdmi_i2c_avalon_slave_0_write),       //                 .write
		.wb_dat_o     (mm_interconnect_1_hdmi_i2c_avalon_slave_0_readdata),    //                 .readdata
		.scl_pad_i    (hdmi_i2c_scl_i),                                        //    conduit_start.scl_i
		.scl_pad_o    (hdmi_i2c_scl_o),                                        //                 .scl_o
		.scl_padoen_o (hdmi_i2c_scl_en),                                       //                 .scl_en
		.sda_pad_i    (hdmi_i2c_sda_i),                                        //                 .sda_i
		.sda_pad_o    (hdmi_i2c_sda_o),                                        //                 .sda_o
		.sda_padoen_o (hdmi_i2c_sda_en),                                       //                 .sda_en
		.wb_inta_o    ()                                                       // interrupt_sender.irq
	);

	MKRVIDOR4000_graphics_lite_sys_irq irq (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_irq_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_irq_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_irq_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_irq_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_irq_s1_readdata),   //                    .readdata
		.in_port    (irq_in_port),                         // external_connection.export
		.out_port   (irq_out_port),                        //                    .export
		.irq        (irq_mapper_receiver1_irq)             //                 irq.irq
	);

	MAILBOX #(
		.pDPRAM_BITS (9),
		.pFIFO_BITS  (4)
	) mb (
		.iCLOCK          (clk_clk),                            //  clock_sink.clk
		.iRESET          (rst_controller_reset_out_reset),     //  reset_sink.reset
		.oMST_AK         (mb_ak),                              // conduit_end.ak
		.iMST_RQ         (mb_rq),                              //            .rq
		.iSLV_WRITE      (mm_interconnect_1_mb_slv_write),     //         slv.write
		.iSLV_READ       (mm_interconnect_1_mb_slv_read),      //            .read
		.iSLV_WRITE_DATA (mm_interconnect_1_mb_slv_writedata), //            .writedata
		.oSLV_READ_DATA  (mm_interconnect_1_mb_slv_readdata),  //            .readdata
		.iSLV_ADDRESS    (mm_interconnect_1_mb_slv_address),   //            .address
		.iMST_WRITE      (mm_interconnect_0_mb_mst_write),     //         mst.write
		.iMST_READ       (mm_interconnect_0_mb_mst_read),      //            .read
		.iMST_WRITE_DATA (mm_interconnect_0_mb_mst_writedata), //            .writedata
		.oMST_READ_DATA  (mm_interconnect_0_mb_mst_readdata),  //            .readdata
		.iMST_ADDRESS    (mm_interconnect_0_mb_mst_address)    //            .address
	);

	tiny_spi #(
		.BAUD_WIDTH (8),
		.BAUD_DIV   (0),
		.SPI_MODE   (0)
	) nina_spi (
		.stb_i (mm_interconnect_1_nina_spi_d_chipselect), //     d.chipselect
		.we_i  (mm_interconnect_1_nina_spi_d_write),      //      .write
		.dat_i (mm_interconnect_1_nina_spi_d_writedata),  //      .writedata
		.adr_i (mm_interconnect_1_nina_spi_d_address),    //      .address
		.dat_o (mm_interconnect_1_nina_spi_d_readdata),   //      .readdata
		.clk_i (clk_clk),                                 //   clk.clk
		.rst_i (rst_controller_reset_out_reset),          // reset.reset
		.int_o (irq_mapper_receiver2_irq),                //   irq.irq
		.MOSI  (nina_spi_MOSI),                           //   spi.MOSI
		.SCLK  (nina_spi_SCLK),                           //      .SCLK
		.MISO  (nina_spi_MISO),                           //      .MISO
		.CS    (nina_spi_CS)                              //      .CS
	);

	MKRVIDOR4000_graphics_lite_sys_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	MKRVIDOR4000_graphics_lite_sys_onchip_memory2_0 onchip_memory2_0 (
		.clk         (clk_clk),                                          //   clk1.clk
		.address     (mm_interconnect_1_onchip_memory2_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_onchip_memory2_0_s1_write),      //       .write
		.readdata    (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),               //       .reset_req
		.address2    (mm_interconnect_1_onchip_memory2_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_1_onchip_memory2_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_1_onchip_memory2_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_1_onchip_memory2_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_1_onchip_memory2_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_1_onchip_memory2_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_1_onchip_memory2_0_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                          //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                   // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	PIO #(
		.pBITS     (32),
		.pMUX_BITS (2)
	) pex_pio (
		.iWRITE      (mm_interconnect_1_pex_pio_s1_write),     //    s1.write
		.iREAD       (mm_interconnect_1_pex_pio_s1_read),      //      .read
		.iWRITE_DATA (mm_interconnect_1_pex_pio_s1_writedata), //      .writedata
		.oREAD_DATA  (mm_interconnect_1_pex_pio_s1_readdata),  //      .readdata
		.iADDRESS    (mm_interconnect_1_pex_pio_s1_address),   //      .address
		.iCLOCK      (clk_clk),                                //   clk.clk
		.iRESET      (rst_controller_reset_out_reset),         // reset.reset
		.iPIO        (pex_pio_in),                             //   pio.in
		.oDIR        (pex_pio_dir),                            //      .dir
		.oPIO        (pex_pio_out),                            //      .out
		.oMUXSEL     (pex_pio_msel)                            //      .msel
	);

	MKRVIDOR4000_graphics_lite_sys_qspi #(
		.DEVICE_FAMILY     ("Cyclone 10 LP"),
		.CS_WIDTH          (3),
		.ADDR_WIDTH        (19),
		.ASI_WIDTH         (4),
		.ASMI_ADDR_WIDTH   (24),
		.ENABLE_4BYTE_ADDR (0),
		.IO_MODE           ("QUAD"),
		.CHIP_SELS         (1),
		.ATOM              ("UNIDIRECTIONAL")
	) qspi (
		.atom_ports_dclk      (qspi_dclk),                                    //       atom_ports.dclk
		.atom_ports_ncs       (qspi_ncs),                                     //                 .ncs
		.atom_ports_oe        (qspi_oe),                                      //                 .oe
		.atom_ports_dataout   (qspi_dataout),                                 //                 .dataout
		.atom_ports_dataoe    (qspi_dataoe),                                  //                 .dataoe
		.atom_ports_datain    (qspi_datain),                                  //                 .datain
		.avl_csr_read         (mm_interconnect_1_qspi_avl_csr_read),          //          avl_csr.read
		.avl_csr_waitrequest  (mm_interconnect_1_qspi_avl_csr_waitrequest),   //                 .waitrequest
		.avl_csr_write        (mm_interconnect_1_qspi_avl_csr_write),         //                 .write
		.avl_csr_addr         (mm_interconnect_1_qspi_avl_csr_address),       //                 .address
		.avl_csr_wrdata       (mm_interconnect_1_qspi_avl_csr_writedata),     //                 .writedata
		.avl_csr_rddata       (mm_interconnect_1_qspi_avl_csr_readdata),      //                 .readdata
		.avl_csr_rddata_valid (mm_interconnect_1_qspi_avl_csr_readdatavalid), //                 .readdatavalid
		.avl_mem_write        (mm_interconnect_1_qspi_avl_mem_write),         //          avl_mem.write
		.avl_mem_burstcount   (mm_interconnect_1_qspi_avl_mem_burstcount),    //                 .burstcount
		.avl_mem_waitrequest  (mm_interconnect_1_qspi_avl_mem_waitrequest),   //                 .waitrequest
		.avl_mem_read         (mm_interconnect_1_qspi_avl_mem_read),          //                 .read
		.avl_mem_addr         (mm_interconnect_1_qspi_avl_mem_address),       //                 .address
		.avl_mem_wrdata       (mm_interconnect_1_qspi_avl_mem_writedata),     //                 .writedata
		.avl_mem_rddata       (mm_interconnect_1_qspi_avl_mem_readdata),      //                 .readdata
		.avl_mem_rddata_valid (mm_interconnect_1_qspi_avl_mem_readdatavalid), //                 .readdatavalid
		.avl_mem_byteenable   (mm_interconnect_1_qspi_avl_mem_byteenable),    //                 .byteenable
		.irq                  (),                                             // interrupt_sender.irq
		.clk                  (clk_0_clk),                                    //       clock_sink.clk
		.reset_n              (~rst_controller_002_reset_out_reset)           //            reset.reset_n
	);

	PIO #(
		.pBITS     (32),
		.pMUX_BITS (2)
	) sam_pio (
		.iWRITE      (mm_interconnect_1_sam_pio_s1_write),     //    s1.write
		.iREAD       (mm_interconnect_1_sam_pio_s1_read),      //      .read
		.iWRITE_DATA (mm_interconnect_1_sam_pio_s1_writedata), //      .writedata
		.oREAD_DATA  (mm_interconnect_1_sam_pio_s1_readdata),  //      .readdata
		.iADDRESS    (mm_interconnect_1_sam_pio_s1_address),   //      .address
		.iCLOCK      (clk_clk),                                //   clk.clk
		.iRESET      (rst_controller_reset_out_reset),         // reset.reset
		.iPIO        (sam_pio_in),                             //   pio.in
		.oDIR        (sam_pio_dir),                            //      .dir
		.oPIO        (sam_pio_out),                            //      .out
		.oMUXSEL     (sam_pio_msel)                            //      .msel
	);

	PWM #(
		.pCHANNELS       (23),
		.pPRESCALER_BITS (32),
		.pMATCH_BITS     (16)
	) sam_pwm (
		.iWRITE_DATA (mm_interconnect_1_sam_pwm_avalon_slave_0_writedata), // avalon_slave_0.writedata
		.iWRITE      (mm_interconnect_1_sam_pwm_avalon_slave_0_write),     //               .write
		.iADDRESS    (mm_interconnect_1_sam_pwm_avalon_slave_0_address),   //               .address
		.iCLOCK      (clk_clk),                                            //     clock_sink.clk
		.iRESET      (rst_controller_reset_out_reset),                     //     reset_sink.reset
		.oPWM        (sam_pwm_pwm)                                         //    conduit_end.pwm
	);

	MKRVIDOR4000_graphics_lite_sys_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_2_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_2_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_2_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_2_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_2_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_2_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_2_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_2_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_2_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	MKRVIDOR4000_graphics_lite_sys_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_0_control_slave_address)   //              .address
	);

	MKRVIDOR4000_graphics_lite_sys_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	PIO #(
		.pBITS     (32),
		.pMUX_BITS (2)
	) wm_pio (
		.iWRITE      (mm_interconnect_1_wm_pio_s1_write),     //    s1.write
		.iREAD       (mm_interconnect_1_wm_pio_s1_read),      //      .read
		.iWRITE_DATA (mm_interconnect_1_wm_pio_s1_writedata), //      .writedata
		.oREAD_DATA  (mm_interconnect_1_wm_pio_s1_readdata),  //      .readdata
		.iADDRESS    (mm_interconnect_1_wm_pio_s1_address),   //      .address
		.iCLOCK      (clk_clk),                               //   clk.clk
		.iRESET      (rst_controller_reset_out_reset),        // reset.reset
		.iPIO        (wm_pio_in),                             //   pio.in
		.oDIR        (wm_pio_dir),                            //      .dir
		.oPIO        (wm_pio_out),                            //      .out
		.oMUXSEL     (wm_pio_msel)                            //      .msel
	);

	MKRVIDOR4000_graphics_lite_sys_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                   (clk_clk),                                 //                                 clk_clk.clk
		.JTAG_BRIDGE_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),          // JTAG_BRIDGE_reset_reset_bridge_in_reset.reset
		.JTAG_BRIDGE_avalon_master_address             (jtag_bridge_avalon_master_address),       //               JTAG_BRIDGE_avalon_master.address
		.JTAG_BRIDGE_avalon_master_waitrequest         (jtag_bridge_avalon_master_waitrequest),   //                                        .waitrequest
		.JTAG_BRIDGE_avalon_master_read                (jtag_bridge_avalon_master_read),          //                                        .read
		.JTAG_BRIDGE_avalon_master_readdata            (jtag_bridge_avalon_master_readdata),      //                                        .readdata
		.JTAG_BRIDGE_avalon_master_readdatavalid       (jtag_bridge_avalon_master_readdatavalid), //                                        .readdatavalid
		.JTAG_BRIDGE_avalon_master_write               (jtag_bridge_avalon_master_write),         //                                        .write
		.JTAG_BRIDGE_avalon_master_writedata           (jtag_bridge_avalon_master_writedata),     //                                        .writedata
		.mb_mst_address                                (mm_interconnect_0_mb_mst_address),        //                                  mb_mst.address
		.mb_mst_write                                  (mm_interconnect_0_mb_mst_write),          //                                        .write
		.mb_mst_read                                   (mm_interconnect_0_mb_mst_read),           //                                        .read
		.mb_mst_readdata                               (mm_interconnect_0_mb_mst_readdata),       //                                        .readdata
		.mb_mst_writedata                              (mm_interconnect_0_mb_mst_writedata)       //                                        .writedata
	);

	MKRVIDOR4000_graphics_lite_sys_mm_interconnect_1 mm_interconnect_1 (
		.clk_clk_clk                                    (clk_clk),                                                    //                                  clk_clk.clk
		.flash_clk_clk_clk                              (clk_0_clk),                                                  //                            flash_clk_clk.clk
		.NEOPIXEL_0_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                             //   NEOPIXEL_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.qspi_reset_reset_bridge_in_reset_reset         (rst_controller_002_reset_out_reset),                         //         qspi_reset_reset_bridge_in_reset.reset
		.NEOPIXEL_0_data_address                        (neopixel_0_data_address),                                    //                          NEOPIXEL_0_data.address
		.NEOPIXEL_0_data_waitrequest                    (neopixel_0_data_waitrequest),                                //                                         .waitrequest
		.NEOPIXEL_0_data_burstcount                     (neopixel_0_data_burstcount),                                 //                                         .burstcount
		.NEOPIXEL_0_data_read                           (neopixel_0_data_read),                                       //                                         .read
		.NEOPIXEL_0_data_readdata                       (neopixel_0_data_readdata),                                   //                                         .readdata
		.NEOPIXEL_0_data_readdatavalid                  (neopixel_0_data_readdatavalid),                              //                                         .readdatavalid
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.csi_i2c_avalon_slave_0_address                 (mm_interconnect_1_csi_i2c_avalon_slave_0_address),           //                   csi_i2c_avalon_slave_0.address
		.csi_i2c_avalon_slave_0_write                   (mm_interconnect_1_csi_i2c_avalon_slave_0_write),             //                                         .write
		.csi_i2c_avalon_slave_0_readdata                (mm_interconnect_1_csi_i2c_avalon_slave_0_readdata),          //                                         .readdata
		.csi_i2c_avalon_slave_0_writedata               (mm_interconnect_1_csi_i2c_avalon_slave_0_writedata),         //                                         .writedata
		.csi_i2c_avalon_slave_0_waitrequest             (~mm_interconnect_1_csi_i2c_avalon_slave_0_waitrequest),      //                                         .waitrequest
		.csi_i2c_avalon_slave_0_chipselect              (mm_interconnect_1_csi_i2c_avalon_slave_0_chipselect),        //                                         .chipselect
		.flash_spi_d_address                            (mm_interconnect_1_flash_spi_d_address),                      //                              flash_spi_d.address
		.flash_spi_d_write                              (mm_interconnect_1_flash_spi_d_write),                        //                                         .write
		.flash_spi_d_readdata                           (mm_interconnect_1_flash_spi_d_readdata),                     //                                         .readdata
		.flash_spi_d_writedata                          (mm_interconnect_1_flash_spi_d_writedata),                    //                                         .writedata
		.flash_spi_d_chipselect                         (mm_interconnect_1_flash_spi_d_chipselect),                   //                                         .chipselect
		.hdmi_i2c_avalon_slave_0_address                (mm_interconnect_1_hdmi_i2c_avalon_slave_0_address),          //                  hdmi_i2c_avalon_slave_0.address
		.hdmi_i2c_avalon_slave_0_write                  (mm_interconnect_1_hdmi_i2c_avalon_slave_0_write),            //                                         .write
		.hdmi_i2c_avalon_slave_0_readdata               (mm_interconnect_1_hdmi_i2c_avalon_slave_0_readdata),         //                                         .readdata
		.hdmi_i2c_avalon_slave_0_writedata              (mm_interconnect_1_hdmi_i2c_avalon_slave_0_writedata),        //                                         .writedata
		.hdmi_i2c_avalon_slave_0_waitrequest            (~mm_interconnect_1_hdmi_i2c_avalon_slave_0_waitrequest),     //                                         .waitrequest
		.hdmi_i2c_avalon_slave_0_chipselect             (mm_interconnect_1_hdmi_i2c_avalon_slave_0_chipselect),       //                                         .chipselect
		.irq_s1_address                                 (mm_interconnect_1_irq_s1_address),                           //                                   irq_s1.address
		.irq_s1_write                                   (mm_interconnect_1_irq_s1_write),                             //                                         .write
		.irq_s1_readdata                                (mm_interconnect_1_irq_s1_readdata),                          //                                         .readdata
		.irq_s1_writedata                               (mm_interconnect_1_irq_s1_writedata),                         //                                         .writedata
		.irq_s1_chipselect                              (mm_interconnect_1_irq_s1_chipselect),                        //                                         .chipselect
		.mb_slv_address                                 (mm_interconnect_1_mb_slv_address),                           //                                   mb_slv.address
		.mb_slv_write                                   (mm_interconnect_1_mb_slv_write),                             //                                         .write
		.mb_slv_read                                    (mm_interconnect_1_mb_slv_read),                              //                                         .read
		.mb_slv_readdata                                (mm_interconnect_1_mb_slv_readdata),                          //                                         .readdata
		.mb_slv_writedata                               (mm_interconnect_1_mb_slv_writedata),                         //                                         .writedata
		.NEOPIXEL_0_csr_address                         (mm_interconnect_1_neopixel_0_csr_address),                   //                           NEOPIXEL_0_csr.address
		.NEOPIXEL_0_csr_write                           (mm_interconnect_1_neopixel_0_csr_write),                     //                                         .write
		.NEOPIXEL_0_csr_read                            (mm_interconnect_1_neopixel_0_csr_read),                      //                                         .read
		.NEOPIXEL_0_csr_readdata                        (mm_interconnect_1_neopixel_0_csr_readdata),                  //                                         .readdata
		.NEOPIXEL_0_csr_writedata                       (mm_interconnect_1_neopixel_0_csr_writedata),                 //                                         .writedata
		.nina_spi_d_address                             (mm_interconnect_1_nina_spi_d_address),                       //                               nina_spi_d.address
		.nina_spi_d_write                               (mm_interconnect_1_nina_spi_d_write),                         //                                         .write
		.nina_spi_d_readdata                            (mm_interconnect_1_nina_spi_d_readdata),                      //                                         .readdata
		.nina_spi_d_writedata                           (mm_interconnect_1_nina_spi_d_writedata),                     //                                         .writedata
		.nina_spi_d_chipselect                          (mm_interconnect_1_nina_spi_d_chipselect),                    //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_1_onchip_memory2_0_s1_address),              //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_1_onchip_memory2_0_s1_write),                //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_1_onchip_memory2_0_s1_readdata),             //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_1_onchip_memory2_0_s1_writedata),            //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_1_onchip_memory2_0_s1_byteenable),           //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_1_onchip_memory2_0_s1_chipselect),           //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_1_onchip_memory2_0_s1_clken),                //                                         .clken
		.onchip_memory2_0_s2_address                    (mm_interconnect_1_onchip_memory2_0_s2_address),              //                      onchip_memory2_0_s2.address
		.onchip_memory2_0_s2_write                      (mm_interconnect_1_onchip_memory2_0_s2_write),                //                                         .write
		.onchip_memory2_0_s2_readdata                   (mm_interconnect_1_onchip_memory2_0_s2_readdata),             //                                         .readdata
		.onchip_memory2_0_s2_writedata                  (mm_interconnect_1_onchip_memory2_0_s2_writedata),            //                                         .writedata
		.onchip_memory2_0_s2_byteenable                 (mm_interconnect_1_onchip_memory2_0_s2_byteenable),           //                                         .byteenable
		.onchip_memory2_0_s2_chipselect                 (mm_interconnect_1_onchip_memory2_0_s2_chipselect),           //                                         .chipselect
		.onchip_memory2_0_s2_clken                      (mm_interconnect_1_onchip_memory2_0_s2_clken),                //                                         .clken
		.pex_pio_s1_address                             (mm_interconnect_1_pex_pio_s1_address),                       //                               pex_pio_s1.address
		.pex_pio_s1_write                               (mm_interconnect_1_pex_pio_s1_write),                         //                                         .write
		.pex_pio_s1_read                                (mm_interconnect_1_pex_pio_s1_read),                          //                                         .read
		.pex_pio_s1_readdata                            (mm_interconnect_1_pex_pio_s1_readdata),                      //                                         .readdata
		.pex_pio_s1_writedata                           (mm_interconnect_1_pex_pio_s1_writedata),                     //                                         .writedata
		.QRCODE_FINDER_0_ctrl_address                   (mm_interconnect_1_qrcode_finder_0_ctrl_address),             //                     QRCODE_FINDER_0_ctrl.address
		.QRCODE_FINDER_0_ctrl_write                     (mm_interconnect_1_qrcode_finder_0_ctrl_write),               //                                         .write
		.QRCODE_FINDER_0_ctrl_read                      (mm_interconnect_1_qrcode_finder_0_ctrl_read),                //                                         .read
		.QRCODE_FINDER_0_ctrl_readdata                  (mm_interconnect_1_qrcode_finder_0_ctrl_readdata),            //                                         .readdata
		.QRCODE_FINDER_0_ctrl_writedata                 (mm_interconnect_1_qrcode_finder_0_ctrl_writedata),           //                                         .writedata
		.qspi_avl_csr_address                           (mm_interconnect_1_qspi_avl_csr_address),                     //                             qspi_avl_csr.address
		.qspi_avl_csr_write                             (mm_interconnect_1_qspi_avl_csr_write),                       //                                         .write
		.qspi_avl_csr_read                              (mm_interconnect_1_qspi_avl_csr_read),                        //                                         .read
		.qspi_avl_csr_readdata                          (mm_interconnect_1_qspi_avl_csr_readdata),                    //                                         .readdata
		.qspi_avl_csr_writedata                         (mm_interconnect_1_qspi_avl_csr_writedata),                   //                                         .writedata
		.qspi_avl_csr_readdatavalid                     (mm_interconnect_1_qspi_avl_csr_readdatavalid),               //                                         .readdatavalid
		.qspi_avl_csr_waitrequest                       (mm_interconnect_1_qspi_avl_csr_waitrequest),                 //                                         .waitrequest
		.qspi_avl_mem_address                           (mm_interconnect_1_qspi_avl_mem_address),                     //                             qspi_avl_mem.address
		.qspi_avl_mem_write                             (mm_interconnect_1_qspi_avl_mem_write),                       //                                         .write
		.qspi_avl_mem_read                              (mm_interconnect_1_qspi_avl_mem_read),                        //                                         .read
		.qspi_avl_mem_readdata                          (mm_interconnect_1_qspi_avl_mem_readdata),                    //                                         .readdata
		.qspi_avl_mem_writedata                         (mm_interconnect_1_qspi_avl_mem_writedata),                   //                                         .writedata
		.qspi_avl_mem_burstcount                        (mm_interconnect_1_qspi_avl_mem_burstcount),                  //                                         .burstcount
		.qspi_avl_mem_byteenable                        (mm_interconnect_1_qspi_avl_mem_byteenable),                  //                                         .byteenable
		.qspi_avl_mem_readdatavalid                     (mm_interconnect_1_qspi_avl_mem_readdatavalid),               //                                         .readdatavalid
		.qspi_avl_mem_waitrequest                       (mm_interconnect_1_qspi_avl_mem_waitrequest),                 //                                         .waitrequest
		.QUAD_ENCODER_0_avalon_slave_0_address          (mm_interconnect_1_quad_encoder_0_avalon_slave_0_address),    //            QUAD_ENCODER_0_avalon_slave_0.address
		.QUAD_ENCODER_0_avalon_slave_0_read             (mm_interconnect_1_quad_encoder_0_avalon_slave_0_read),       //                                         .read
		.QUAD_ENCODER_0_avalon_slave_0_readdata         (mm_interconnect_1_quad_encoder_0_avalon_slave_0_readdata),   //                                         .readdata
		.sam_pio_s1_address                             (mm_interconnect_1_sam_pio_s1_address),                       //                               sam_pio_s1.address
		.sam_pio_s1_write                               (mm_interconnect_1_sam_pio_s1_write),                         //                                         .write
		.sam_pio_s1_read                                (mm_interconnect_1_sam_pio_s1_read),                          //                                         .read
		.sam_pio_s1_readdata                            (mm_interconnect_1_sam_pio_s1_readdata),                      //                                         .readdata
		.sam_pio_s1_writedata                           (mm_interconnect_1_sam_pio_s1_writedata),                     //                                         .writedata
		.sam_pwm_avalon_slave_0_address                 (mm_interconnect_1_sam_pwm_avalon_slave_0_address),           //                   sam_pwm_avalon_slave_0.address
		.sam_pwm_avalon_slave_0_write                   (mm_interconnect_1_sam_pwm_avalon_slave_0_write),             //                                         .write
		.sam_pwm_avalon_slave_0_writedata               (mm_interconnect_1_sam_pwm_avalon_slave_0_writedata),         //                                         .writedata
		.SDRAM_ARBITER_avl_address                      (mm_interconnect_1_sdram_arbiter_avl_address),                //                        SDRAM_ARBITER_avl.address
		.SDRAM_ARBITER_avl_write                        (mm_interconnect_1_sdram_arbiter_avl_write),                  //                                         .write
		.SDRAM_ARBITER_avl_read                         (mm_interconnect_1_sdram_arbiter_avl_read),                   //                                         .read
		.SDRAM_ARBITER_avl_readdata                     (mm_interconnect_1_sdram_arbiter_avl_readdata),               //                                         .readdata
		.SDRAM_ARBITER_avl_writedata                    (mm_interconnect_1_sdram_arbiter_avl_writedata),              //                                         .writedata
		.SDRAM_ARBITER_avl_burstcount                   (mm_interconnect_1_sdram_arbiter_avl_burstcount),             //                                         .burstcount
		.SDRAM_ARBITER_avl_byteenable                   (mm_interconnect_1_sdram_arbiter_avl_byteenable),             //                                         .byteenable
		.SDRAM_ARBITER_avl_readdatavalid                (mm_interconnect_1_sdram_arbiter_avl_readdatavalid),          //                                         .readdatavalid
		.SDRAM_ARBITER_avl_waitrequest                  (mm_interconnect_1_sdram_arbiter_avl_waitrequest),            //                                         .waitrequest
		.sysid_qsys_0_control_slave_address             (mm_interconnect_1_sysid_qsys_0_control_slave_address),       //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_1_sysid_qsys_0_control_slave_readdata),      //                                         .readdata
		.timer_0_s1_address                             (mm_interconnect_1_timer_0_s1_address),                       //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_1_timer_0_s1_write),                         //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_1_timer_0_s1_readdata),                      //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_1_timer_0_s1_writedata),                     //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_1_timer_0_s1_chipselect),                    //                                         .chipselect
		.wm_pio_s1_address                              (mm_interconnect_1_wm_pio_s1_address),                        //                                wm_pio_s1.address
		.wm_pio_s1_write                                (mm_interconnect_1_wm_pio_s1_write),                          //                                         .write
		.wm_pio_s1_read                                 (mm_interconnect_1_wm_pio_s1_read),                           //                                         .read
		.wm_pio_s1_readdata                             (mm_interconnect_1_wm_pio_s1_readdata),                       //                                         .readdata
		.wm_pio_s1_writedata                            (mm_interconnect_1_wm_pio_s1_writedata)                       //                                         .writedata
	);

	MKRVIDOR4000_graphics_lite_sys_mm_interconnect_2 mm_interconnect_2 (
		.clk_clk_clk                                     (clk_clk),                                  //                                   clk_clk.clk
		.SDRAM_ARBITER_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),           // SDRAM_ARBITER_reset_reset_bridge_in_reset.reset
		.SDRAM_ARBITER_sdram_address                     (sdram_arbiter_sdram_address),              //                       SDRAM_ARBITER_sdram.address
		.SDRAM_ARBITER_sdram_waitrequest                 (sdram_arbiter_sdram_waitrequest),          //                                          .waitrequest
		.SDRAM_ARBITER_sdram_byteenable                  (sdram_arbiter_sdram_byteenable),           //                                          .byteenable
		.SDRAM_ARBITER_sdram_read                        (sdram_arbiter_sdram_read),                 //                                          .read
		.SDRAM_ARBITER_sdram_readdata                    (sdram_arbiter_sdram_readdata),             //                                          .readdata
		.SDRAM_ARBITER_sdram_readdatavalid               (sdram_arbiter_sdram_readdatavalid),        //                                          .readdatavalid
		.SDRAM_ARBITER_sdram_write                       (sdram_arbiter_sdram_write),                //                                          .write
		.SDRAM_ARBITER_sdram_writedata                   (sdram_arbiter_sdram_writedata),            //                                          .writedata
		.sdram_s1_address                                (mm_interconnect_2_sdram_s1_address),       //                                  sdram_s1.address
		.sdram_s1_write                                  (mm_interconnect_2_sdram_s1_write),         //                                          .write
		.sdram_s1_read                                   (mm_interconnect_2_sdram_s1_read),          //                                          .read
		.sdram_s1_readdata                               (mm_interconnect_2_sdram_s1_readdata),      //                                          .readdata
		.sdram_s1_writedata                              (mm_interconnect_2_sdram_s1_writedata),     //                                          .writedata
		.sdram_s1_byteenable                             (mm_interconnect_2_sdram_s1_byteenable),    //                                          .byteenable
		.sdram_s1_readdatavalid                          (mm_interconnect_2_sdram_s1_readdatavalid), //                                          .readdatavalid
		.sdram_s1_waitrequest                            (mm_interconnect_2_sdram_s1_waitrequest),   //                                          .waitrequest
		.sdram_s1_chipselect                             (mm_interconnect_2_sdram_s1_chipselect)     //                                          .chipselect
	);

	MKRVIDOR4000_graphics_lite_sys_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_0_clk),                          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule

// forearm_control.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module forearm_control (
		input  wire        clk_clk,                                       //                         clk.clk
		input  wire [15:0] myocontrol_0_avalon_slave_0_address,           // myocontrol_0_avalon_slave_0.address
		input  wire        myocontrol_0_avalon_slave_0_write,             //                            .write
		input  wire [31:0] myocontrol_0_avalon_slave_0_writedata,         //                            .writedata
		input  wire        myocontrol_0_avalon_slave_0_read,              //                            .read
		output wire [31:0] myocontrol_0_avalon_slave_0_readdata,          //                            .readdata
		output wire        myocontrol_0_avalon_slave_0_waitrequest,       //                            .waitrequest
		input  wire        myocontrol_0_conduit_end_angle_miso,           //    myocontrol_0_conduit_end.angle_miso
		output wire        myocontrol_0_conduit_end_angle_mosi,           //                            .angle_mosi
		output wire        myocontrol_0_conduit_end_angle_sck,            //                            .angle_sck
		output wire [2:0]  myocontrol_0_conduit_end_angle_ss_n_o,         //                            .angle_ss_n_o
		output wire        myocontrol_0_conduit_end_gpio_n,               //                            .gpio_n
		input  wire        myocontrol_0_conduit_end_mirrored_muscle_unit, //                            .mirrored_muscle_unit
		input  wire        myocontrol_0_conduit_end_miso,                 //                            .miso
		output wire        myocontrol_0_conduit_end_mosi,                 //                            .mosi
		input  wire        myocontrol_0_conduit_end_power_sense_n,        //                            .power_sense_n
		output wire [2:0]  myocontrol_0_conduit_end_ss_n_o,               //                            .ss_n_o
		output wire        myocontrol_0_conduit_end_sck,                  //                            .sck
		input  wire        reset_reset_n                                  //                       reset.reset_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> MYOControl_0:reset

	MYOControl #(
		.NUMBER_OF_MOTORS        (3),
		.CLOCK_SPEED_HZ          (48000000),
		.ENABLE_MYOBRICK_CONTROL (0)
	) myocontrol_0 (
		.reset                (rst_controller_reset_out_reset),                //          reset.reset
		.address              (myocontrol_0_avalon_slave_0_address),           // avalon_slave_0.address
		.write                (myocontrol_0_avalon_slave_0_write),             //               .write
		.writedata            (myocontrol_0_avalon_slave_0_writedata),         //               .writedata
		.read                 (myocontrol_0_avalon_slave_0_read),              //               .read
		.readdata             (myocontrol_0_avalon_slave_0_readdata),          //               .readdata
		.waitrequest          (myocontrol_0_avalon_slave_0_waitrequest),       //               .waitrequest
		.angle_miso           (myocontrol_0_conduit_end_angle_miso),           //    conduit_end.angle_miso
		.angle_mosi           (myocontrol_0_conduit_end_angle_mosi),           //               .angle_mosi
		.angle_sck            (myocontrol_0_conduit_end_angle_sck),            //               .angle_sck
		.angle_ss_n_o         (myocontrol_0_conduit_end_angle_ss_n_o),         //               .angle_ss_n_o
		.gpio_n               (myocontrol_0_conduit_end_gpio_n),               //               .gpio_n
		.mirrored_muscle_unit (myocontrol_0_conduit_end_mirrored_muscle_unit), //               .mirrored_muscle_unit
		.miso                 (myocontrol_0_conduit_end_miso),                 //               .miso
		.mosi                 (myocontrol_0_conduit_end_mosi),                 //               .mosi
		.power_sense_n        (myocontrol_0_conduit_end_power_sense_n),        //               .power_sense_n
		.ss_n_o               (myocontrol_0_conduit_end_ss_n_o),               //               .ss_n_o
		.sck                  (myocontrol_0_conduit_end_sck),                  //               .sck
		.clock                (clk_clk)                                        //     clock_sink.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule

// MKRVIDOR4000_mipi.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module MKRVIDOR4000_mipi (
		input  wire        arb_fb_clk,     //   arb_fb.clk
		input  wire        arb_fb_rdy,     //         .rdy
		output wire [30:0] arb_fb_data,    //         .data
		output wire        arb_fb_dv,      //         .dv
		output wire        arb_fb_start,   //         .start
		input  wire        arb_mipi_clk,   // arb_mipi.clk
		input  wire [14:0] arb_mipi_data,  //         .data
		input  wire        arb_mipi_dv,    //         .dv
		input  wire        arb_mipi_start, //         .start
		input  wire        clk_clk,        //      clk.clk
		input  wire        fb_st_start,    //    fb_st.start
		input  wire [30:0] fb_st_data,     //         .data
		input  wire        fb_st_dv,       //         .dv
		output wire        fb_st_ready,    //         .ready
		output wire [7:0]  fb_vport_blu,   // fb_vport.blu
		output wire        fb_vport_de,    //         .de
		output wire [7:0]  fb_vport_grn,   //         .grn
		output wire        fb_vport_hs,    //         .hs
		output wire        fb_vport_vs,    //         .vs
		output wire [7:0]  fb_vport_red,   //         .red
		input  wire        mipi_rx_clk,    //  mipi_rx.clk
		input  wire [1:0]  mipi_rx_data,   //         .data
		output wire [23:0] mipi_st_data,   //  mipi_st.data
		output wire        mipi_st_start,  //         .start
		output wire        mipi_st_dv,     //         .dv
		input  wire        reset_reset_n,  //    reset.reset_n
		output wire [11:0] sdram_addr,     //    sdram.addr
		output wire [1:0]  sdram_ba,       //         .ba
		output wire        sdram_cas_n,    //         .cas_n
		output wire        sdram_cke,      //         .cke
		output wire        sdram_cs_n,     //         .cs_n
		inout  wire [15:0] sdram_dq,       //         .dq
		output wire [1:0]  sdram_dqm,      //         .dqm
		output wire        sdram_ras_n,    //         .ras_n
		output wire        sdram_we_n,     //         .we_n
		input  wire        vid_clk         //      vid.clk
	);

	wire  [15:0] sdram_arbiter_sdram_readdata;             // mm_interconnect_0:SDRAM_ARBITER_sdram_readdata -> SDRAM_ARBITER:iSDRAM_READ_DATA
	wire         sdram_arbiter_sdram_waitrequest;          // mm_interconnect_0:SDRAM_ARBITER_sdram_waitrequest -> SDRAM_ARBITER:iSDRAM_WAIT_REQUEST
	wire  [21:0] sdram_arbiter_sdram_address;              // SDRAM_ARBITER:oSDRAM_ADDRESS -> mm_interconnect_0:SDRAM_ARBITER_sdram_address
	wire         sdram_arbiter_sdram_read;                 // SDRAM_ARBITER:oSDRAM_READ -> mm_interconnect_0:SDRAM_ARBITER_sdram_read
	wire   [1:0] sdram_arbiter_sdram_byteenable;           // SDRAM_ARBITER:oSDRAM_BYTE_ENABLE -> mm_interconnect_0:SDRAM_ARBITER_sdram_byteenable
	wire         sdram_arbiter_sdram_readdatavalid;        // mm_interconnect_0:SDRAM_ARBITER_sdram_readdatavalid -> SDRAM_ARBITER:iSDRAM_READ_DATA_VALID
	wire         sdram_arbiter_sdram_write;                // SDRAM_ARBITER:oSDRAM_WRITE -> mm_interconnect_0:SDRAM_ARBITER_sdram_write
	wire  [15:0] sdram_arbiter_sdram_writedata;            // SDRAM_ARBITER:oSDRAM_WRITE_DATA -> mm_interconnect_0:SDRAM_ARBITER_sdram_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;    // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;      // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;   // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;       // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;          // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;    // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid; // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;         // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;     // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         rst_controller_reset_out_reset;           // rst_controller:reset_out -> [SDRAM_ARBITER:iRESET, mm_interconnect_0:SDRAM_ARBITER_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	FBST #(
		.pHRES   (640),
		.pVRES   (480),
		.pHTOTAL (762),
		.pVTOTAL (525),
		.pHSS    (656),
		.pHSE    (752),
		.pVSS    (490),
		.pVSE    (492)
	) fbst_0 (
		.oBLU          (fb_vport_blu), //   vport.blu
		.oDE           (fb_vport_de),  //        .de
		.oGRN          (fb_vport_grn), //        .grn
		.oHS           (fb_vport_hs),  //        .hs
		.oVS           (fb_vport_vs),  //        .vs
		.oRED          (fb_vport_red), //        .red
		.iCLK          (vid_clk),      // vid_clk.clk
		.iFB_START     (fb_st_start),  //  stream.start
		.iFB_DATA      (fb_st_data),   //        .data
		.iFB_DATAVALID (fb_st_dv),     //        .dv
		.oFB_READY     (fb_st_ready)   //        .ready
	);

	MIPI_RX mipi_rx_st_0 (
		.iMIPI_CLK       (mipi_rx_clk),   //    mipi.clk
		.iMIPI_D         (mipi_rx_data),  //        .data
		.oMIPI_DATA      (mipi_st_data),  // mipi_st.data
		.oMIPI_START     (mipi_st_start), //        .start
		.oMIPI_DATAVALID (mipi_st_dv)     //        .dv
	);

	SDRAM_ARBITER #(
		.pBURST_SIZE   (128),
		.pCAM_OFFSET_A (0),
		.pCAM_OFFSET_B (307200),
		.pFB_OFFSET    (614400),
		.pFB_SIZE      (307200),
		.pADDRESS_BITS (22)
	) sdram_arbiter (
		.oSDRAM_ADDRESS         (sdram_arbiter_sdram_address),       // sdram.address
		.oSDRAM_WRITE           (sdram_arbiter_sdram_write),         //      .write
		.oSDRAM_READ            (sdram_arbiter_sdram_read),          //      .read
		.oSDRAM_WRITE_DATA      (sdram_arbiter_sdram_writedata),     //      .writedata
		.iSDRAM_READ_DATA       (sdram_arbiter_sdram_readdata),      //      .readdata
		.iSDRAM_WAIT_REQUEST    (sdram_arbiter_sdram_waitrequest),   //      .waitrequest
		.iSDRAM_READ_DATA_VALID (sdram_arbiter_sdram_readdatavalid), //      .readdatavalid
		.oSDRAM_BYTE_ENABLE     (sdram_arbiter_sdram_byteenable),    //      .byteenable
		.iMEM_CLK               (clk_clk),                           // clock.clk
		.iRESET                 (rst_controller_reset_out_reset),    // reset.reset
		.iFB_CLK                (arb_fb_clk),                        //    fb.clk
		.iFB_READY              (arb_fb_rdy),                        //      .rdy
		.oFB_DATA               (arb_fb_data),                       //      .data
		.oFB_DATA_VALID         (arb_fb_dv),                         //      .dv
		.oFB_START              (arb_fb_start),                      //      .start
		.iMIPI_CLK              (arb_mipi_clk),                      //  mipi.clk
		.iMIPI_DATA             (arb_mipi_data),                     //      .data
		.iMIPI_DATA_VALID       (arb_mipi_dv),                       //      .dv
		.iMIPI_START            (arb_mipi_start),                    //      .start
		.oAVL_READ_DATA         (),                                  //   avl.readdata
		.oAVL_READ_DATA_VALID   (),                                  //      .readdatavalid
		.iAVL_WRITE_DATA        (),                                  //      .writedata
		.oAVL_WAIT_REQUEST      (),                                  //      .waitrequest
		.iAVL_ADDRESS           (),                                  //      .address
		.iAVL_BURST_COUNT       (),                                  //      .burstcount
		.iAVL_READ              (),                                  //      .read
		.iAVL_WRITE             (),                                  //      .write
		.iAVL_BYTE_ENABLE       ()                                   //      .byteenable
	);

	MKRVIDOR4000_mipi_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	MKRVIDOR4000_mipi_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                     (clk_clk),                                  //                                   clk_clk.clk
		.SDRAM_ARBITER_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),           // SDRAM_ARBITER_reset_reset_bridge_in_reset.reset
		.SDRAM_ARBITER_sdram_address                     (sdram_arbiter_sdram_address),              //                       SDRAM_ARBITER_sdram.address
		.SDRAM_ARBITER_sdram_waitrequest                 (sdram_arbiter_sdram_waitrequest),          //                                          .waitrequest
		.SDRAM_ARBITER_sdram_byteenable                  (sdram_arbiter_sdram_byteenable),           //                                          .byteenable
		.SDRAM_ARBITER_sdram_read                        (sdram_arbiter_sdram_read),                 //                                          .read
		.SDRAM_ARBITER_sdram_readdata                    (sdram_arbiter_sdram_readdata),             //                                          .readdata
		.SDRAM_ARBITER_sdram_readdatavalid               (sdram_arbiter_sdram_readdatavalid),        //                                          .readdatavalid
		.SDRAM_ARBITER_sdram_write                       (sdram_arbiter_sdram_write),                //                                          .write
		.SDRAM_ARBITER_sdram_writedata                   (sdram_arbiter_sdram_writedata),            //                                          .writedata
		.sdram_s1_address                                (mm_interconnect_0_sdram_s1_address),       //                                  sdram_s1.address
		.sdram_s1_write                                  (mm_interconnect_0_sdram_s1_write),         //                                          .write
		.sdram_s1_read                                   (mm_interconnect_0_sdram_s1_read),          //                                          .read
		.sdram_s1_readdata                               (mm_interconnect_0_sdram_s1_readdata),      //                                          .readdata
		.sdram_s1_writedata                              (mm_interconnect_0_sdram_s1_writedata),     //                                          .writedata
		.sdram_s1_byteenable                             (mm_interconnect_0_sdram_s1_byteenable),    //                                          .byteenable
		.sdram_s1_readdatavalid                          (mm_interconnect_0_sdram_s1_readdatavalid), //                                          .readdatavalid
		.sdram_s1_waitrequest                            (mm_interconnect_0_sdram_s1_waitrequest),   //                                          .waitrequest
		.sdram_s1_chipselect                             (mm_interconnect_0_sdram_s1_chipselect)     //                                          .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
